`define OPCODE_WIDTH 6
`define RTYPE 6'h0
`define BEQ 6'h4
`define BNE 6'h5
`define ORI 6'hd
`define LUI 6'hf
`define JAL 6'h3
`define SLTI 6'ha
`define ADDI 6'h8
`define ANDI 6'hc
`define ADDIU 6'h9
`define SLTIU 6'hb
`define STORE_WORD 6'h2b
`define STORE_BYTE 6'h2c
`define STORE_HALF 6'h2d
`define LOAD_WORD 6'h23
`define LOAD_BYTE 6'h26
`define LOAD_HALF 6'h27
`define LOAD_BYTE_UNSIGNED 6'h24
`define LOAD_HALF_UNSIGNED 6'h25

`define FUNCT_WIDTH 6
`define ADD 6'b100000
`define SUB 6'b100010
`define SUBU 6'b100011
`define AND 6'b100100
`define OR 6'b100101
`define NOR 6'b100111
`define SLT 6'b101010
`define SLTU 6'b101011
`define SLL 6'b000000
`define SRL 6'b000010
`define SRA 6'b101001
`define EQ 6'b001100
`define NEQ 6'b001101
`define GE 6'b101100
`define GEU 6'b101101
`define ADDU 6'b100001
`define JR 6'b001000

`define DWIDTH 32
`define IWIDTH 32
`define AWIDTH 5
`define PC_WIDTH 32
`define AWIDTH_MEM 32
`define IMM_WIDTH 16
`define ALU_CONTROL 5
`define JUMP_WIDTH 26
`define DEPTH 4